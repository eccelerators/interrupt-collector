-- ******************************************************************************
-- 
--                   /------o
--             eccelerators
--          o------/
-- 
--  This file is an Eccelerators GmbH sample project.
-- 
--  MIT License:
--  Copyright (c) 2023 Eccelerators GmbH
-- 
--  Permission is hereby granted, free of charge, to any person obtaining a copy
--  of this software and associated documentation files (the "Software"), to deal
--  in the Software without restriction, including without limitation the rights
--  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
--  copies of the Software, and to permit persons to whom the Software is
--  furnished to do so, subject to the following conditions:
-- 
--  The above copyright notice and this permission notice shall be included in all
--  copies or substantial portions of the Software.
-- 
--  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
--  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
--  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
--  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
--  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
--  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
--  SOFTWARE.
-- ******************************************************************************
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    
use work.EventCatcherIfcPackage.all;
use work.tb_bus_pkg.all;
use work.tb_signals_pkg.all;
use work.tb_base_pkg.all;


entity tb_top_wishbone is
    generic (
        stimulus_path : string := "../../tb/simstm/";
        stimulus_file : string := "TestMainWishbone.stm"
    );
end;

architecture behavioural of tb_top_wishbone is

    signal simdone : std_logic := '0';
    
    signal Clk : std_logic := '0';
    signal Rst : std_logic := '1';
    signal TimeoutAck_Detected : std_logic := '0';
    signal TimeoutAck_Rec_Clear : std_logic := '0';
    
    signal executing_line : integer := 0;
    signal executing_file : text_line;
    signal marker : std_logic_vector(15 downto 0) := (others => '0');
    
    signal signals_in : t_signals_in;
    signal signals_out : t_signals_out;

    signal bus_down : t_bus_down;
    signal bus_up : t_bus_up;    
    
    signal EventCatcherIfcWishboneDown : T_EventCatcherIfcWishboneDown;
    signal EventCatcherIfcWishboneUp : T_EventCatcherIfcWishboneUp;    
    
    signal EventCatcherIfcEventCatcherBlkDown :T_EventCatcherIfcEventCatcherBlkDown;
    signal EventCatcherIfcEventCatcherBlkUp : T_EventCatcherIfcEventCatcherBlkUp;
    signal EventCatcherIfcTrace : T_EventCatcherIfcTrace;
    
    signal EventOut : std_logic_vector(3 downto 0);
    signal PreviousEventOut0 : std_logic;
    signal EventCatch : std_logic_vector(3 downto 0);
    signal EventPuls : std_logic_vector(3 downto 0);
    signal EventPuls0 : std_logic;
    signal EventPuls1 : std_logic;
    signal EventPuls2 : std_logic;
    signal EventPuls3 : std_logic;
    
begin

    Rst <= transport '0' after 100 ns;
    Clk <= transport (not Clk) and (not SimDone)  after 10 ns / 2; -- 100MHz
    
    EventOut <= signals_out.EventOut_4;

    signals_in.in_signal <= '0';
    signals_in.in_signal_1 <= (others => '0');
    signals_in.in_signal_2 <= '0';
    signals_in.in_signal_3 <= '0';
    signals_in.EventCatch_4 <= EventCatch;
    
    EventPuls <= EventPuls3 & EventPuls2 & EventPuls1 & EventPuls0;
    
    EventPuls1 <= EventPuls0 or (EventOut(1) and EventCatcherIfcEventCatcherBlkDown.WTransPulseEventCatchReg); --generate event at same clock as event confirm
    
    
    EventPuls3 <= EventPuls0 or (EventOut(3) and EventCatcherIfcEventCatcherBlkDown.WTransPulseEventOverrunReg); --generate event at same clock as overrun confirm
    
    
    prcGenEventPulses : process ( Clk, Rst) is
    begin
        if Rst then
        
            EventPuls0 <= '0';
            EventPuls2 <= '0';
            PreviousEventOut0 <= '0';
            
        elsif rising_edge(Clk) then
        
            PreviousEventOut0 <= EventOut(0);
            EventPuls0 <= '0'; -- default assignment
            EventPuls2 <= '0'; -- default assignment
            
            if not PreviousEventOut0 and EventOut(0) then
                EventPuls0 <= '1'; --generate event at all at rising EventOut0 edge
            end if;
            
            if EventCatcherIfcEventCatcherBlkDown.WTransPulseEventCatchReg and EventOut(2) then
                EventPuls2 <= '1'; 
            end if; --generate event one clock after event confirm
            
        end if;  
    end process;
    
    i_tb_simstm : entity work.tb_simstm
        generic map (
            stimulus_path => stimulus_path,
            stimulus_file => stimulus_file          
        )
        port map (
            clk => Clk,
            rst => Rst,
            simdone => SimDone,       
            executing_line => executing_line,
            executing_file => executing_file,
            marker => marker,
            signals_in => signals_in,
            signals_out => signals_out,
            bus_down => bus_down,
            bus_up => bus_up
        );
        
    EventCatcherIfcWishboneDown.Adr <= bus_down.wishbone.adr(EventCatcherIfcWishboneDown.Adr'LENGTH - 1 downto 0);
    EventCatcherIfcWishboneDown.Sel <= bus_down.wishbone.sel;
    EventCatcherIfcWishboneDown.DatIn <= bus_down.wishbone.data;
    EventCatcherIfcWishboneDown.We <= bus_down.wishbone.we;
    EventCatcherIfcWishboneDown.Stb <= bus_down.wishbone.stb;
    EventCatcherIfcWishboneDown.Cyc <= bus_down.wishbone.cyc;
    
    bus_up.wishbone.data <= EventCatcherIfcWishboneUp.DatOut;
    bus_up.wishbone.ack <= EventCatcherIfcWishboneUp.Ack;
    
    
    i_EventCatcherIfcWishbone : entity work.EventCatcherIfcWishbone
        port map(
            Clk => Clk,
            Rst => Rst,
            WishboneDown => EventCatcherIfcWishboneDown,
            WishboneUp => EventCatcherIfcWishboneUp,
            Trace => EventCatcherIfcTrace,
            EventCatcherBlkDown => EventCatcherIfcEventCatcherBlkDown,
            EventCatcherBlkUp => EventCatcherIfcEventCatcherBlkUp
        );

                    
    i_EventCatcher: entity work.EventCatcher
    generic map (
        BIT_WIDTH => 4
    )
    port map(
        Clk => Clk,
        Rst => Rst,
        EventPuls => EventPuls,
        EventCatch => EventCatch,
        Mask => EventCatcherIfcEventCatcherBlkDown.Mask,
        CatchWritten => EventCatcherIfcEventCatcherBlkDown.CatchWritten,
        WTransPulseEventCatchReg => EventCatcherIfcEventCatcherBlkDown.WTransPulseEventCatchReg,
        CatchToBeRead => EventCatcherIfcEventCatcherBlkUp.CatchToBeRead,
        OverrunWritten => EventCatcherIfcEventCatcherBlkDown.OverrunWritten,
        WTransPulseEventOverrunReg => EventCatcherIfcEventCatcherBlkDown.WTransPulseEventOverrunReg,
        OverrunToBeRead => EventCatcherIfcEventCatcherBlkUp.OverrunToBeRead
    );
  
end;